// you're a senior FPGA Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Create 8 D flip-flops with active high synchronous reset. The flip-flops must be reset to 0x34 rather than zero. All DFFs should be triggered by the negative edge of clk.

// Hint: Resetting a register to '1' is sometimes called "preset"

module top_module (
    input clk,
    input reset,
    input [7:0] d,
    output [7:0] q
);

	// Insert your code here

endmodule
