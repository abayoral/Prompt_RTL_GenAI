// you're a senior FPGA Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Make 3 instances of full-adder to create a 3-bit binary ripple-carry adder. 
// The adder adds two 3-bit numbers and a carry-in to produce a 3-bit sum and carry out. 
// To encourage you to actually instantiate full adders, also output the carry-out from 
// each full adder in the ripple-carry adder. cout[2] is the final carry-out from the last 
// full adder, and is the carry-out you usually see.

module top_module( 
    input [2:0] a, b,
    input cin,
    output [2:0] cout,
    output [2:0] sum );

    // Insert your code here

endmodule


