// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Create a module with 3 inputs and 4 outputs that behaves like wires that makes these connections:

// a -> w
// b -> x
// b -> y
// c -> z

// Hint: The concatenation operator { signal1, signal2, signal3, ... } would be useful here.

module top_module( 
    input a,b,c,
    output w,x,y,z );

// Insert your code here

endmodule
