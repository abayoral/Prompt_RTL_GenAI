// Imagine you hold the position of a senior Digital Design Engineer at a leading hardware design company, and you are entrusted with the mission of creating a crucial module in Verilog for an upcoming product that is key to the future of your company's esteemed position within the computer hardware industry. The functionality and reliability of this module are paramount, as it will directly affect the company's standing and credibility in a highly competitive market.

// Your task involves designing a group of 8 D flip-flops (DFFs), each with an active high synchronous reset feature. The D flip-flops should all be activated by the positive edge of the clock signal (clk), meaning they will capture the input data at the rising edge of each clock cycle. The synchronous reset implies that the reset condition will only take effect on the active edge of the clock, ensuring proper timing and control within your digital design system.

// Specifically, you are expected to complete the Verilog module outlined below, where the module is named `top_module`. It takes an 8-bit input vector `d`, a clock input `clk`, and a reset input `reset`, and it should produce an 8-bit output vector `q` that reflects the stored state of each corresponding D flip-flop. It is up to you to decide how best to implement this functionality within the given code structure.

// module top_module (
//     input clk,
//     input reset,            // Synchronous reset
//     input [7:0] d,
//     output [7:0] q
// );

// Insert your code here

// endmodule