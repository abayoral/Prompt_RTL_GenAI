module top_module(
    input clk,
    input [7:0] in,
    input reset,    // Synchronous reset
    output reg [23:0] out_bytes,
    output reg done); //

    // State enumeration
    typedef enum reg [1:0] {
        IDLE = 2'b00,
        BYTE1 = 2'b01,
        BYTE2 = 2'b10,
        BYTE3 = 2'b11
    } state_t;
    
    state_t state, next_state;
    reg [23:0] message_reg;
    
    // State transition logic (FSM)
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            state <= IDLE;
        end
        else begin
            state <= next_state;
        end
    end

    // Next state and output logic
    always @(*) begin
        // Default values
        done = 0;
        next_state = state;
        
        case (state)
            IDLE: begin
                if (in[3] == 1) begin
                    next_state = BYTE1;
                end
            end
            BYTE1: begin
                next_state = BYTE2;
            end
            BYTE2: begin
                next_state = BYTE3;
            end
            BYTE3: begin
                next_state = IDLE;
                done = 1;
            end
        endcase
    end

    // Datapath to accumulate bytes
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            message_reg <= 24'b0;
            out_bytes <= 24'b0;
        end
        else begin
            case (next_state)
                IDLE: begin
                    // Clear message register in IDLE state
                    message_reg <= 24'b0;
                end
                BYTE1: begin
                    message_reg[23:16] <= in;
                end
                BYTE2: begin
                    message_reg[15:8] <= in;
                end
                BYTE3: begin
                    message_reg[7:0] <= in;
                    out_bytes <= {message_reg[23:8], in};
                end
            endcase

            if (done) begin
                out_bytes <= message_reg;
            end
        end
    end
endmodule