Imagine you are a highly experienced Digital Logic Design Engineer at a top-tier hardware design firm. Your current assignment involves designing a critical Verilog module that will be integral to a next-generation computer hardware product. The module's successful performance is crucial, as it will greatly influence the company's standing in the industry.

The specific task is centered on creating a "population count" circuit—a type of combinational logic design that determines how many bits in a binary vector are set to '1'. In this case, your circuit will need to evaluate a 3-bit input vector. Based on the number of bits that are '1', the circuit should produce an output. 

Your Verilog module, named top_module, is defined with a 3-bit input vector (in) and a 2-bit output vector (out). Within this module, you will need to insert your design logic where indicated. Although the problem statement is concise, keep in mind that your implementation must accurately count the number of '1's in the provided 3-bit input and output the result as a 2-bit binary number.

Your expanded assignment is as follows:

• As a lead engineer, your goal is to implement and validate a population count circuit using Verilog.  
• The circuit should accept a 3-bit input vector labeled "in".  
• It must calculate the count of bits set to '1' within this input.  
• The resulting count, represented as a 2-bit binary value, should be output via the "out" port.  
• Begin your module definition with the provided top_module template, and integrate your solution where the comment "INSERT YOUR CODE HERE" is indicated.

This task challenges you to apply your logic design expertise to ensure the module is both efficient and reliable for its intended application. No additional functionality or extraneous outputs are necessary beyond the proper counting of '1' bits and mapping that count to a 2-bit output.