Imagine you are a senior Digital Design Engineer at a prominent hardware design company, and one of your key responsibilities is to create an essential Verilog module for an upcoming, cutting-edge product. The delivery and performance of this module are crucial to maintaining your company’s esteemed status within the competitive computer hardware sector.

The module you are tasked to develop involves interaction with the PS/2 mouse protocol, which is known to transmit data in messages of precisely three bytes. Within the continuous stream of incoming bytes, it’s not inherently clear where a specific message begins or ends. The only distinguishing factor is that the first byte of each three-byte message consistently has bit[3]=1. For the subsequent two bytes of the message, bit[3] can either be 1 or 0, as this depends on the actual data being transmitted.

The goal is to design a finite state machine (FSM) that will scrutinize this byte stream and accurately identify message boundaries. The method you’ll use involves disregarding bytes until a byte with bit[3]=1 is detected. Upon sensing such a byte, it is presumed to be the initial byte of a new message, and a signal is emitted indicating the completion of receiving a message once all three bytes have been successfully captured.

Building upon the existing state machine that effectively discerns three-byte messages within the PS/2 byte stream, the next step is to enhance this framework by incorporating a datapath. This additional functionality will enable the module to output the entire 24-bit message (comprised of the 3 bytes) once a packet is fully received. Here, the output should be structured such that out_bytes[23:16] represents the first byte, out_bytes[15:8] encapsulates the second byte, and out_bytes[7:0] stores the final byte.

It's important to note that the output out_bytes must be valid and convey the complete message precisely at the moment when the done signal is asserted. At other times, what is outputted is not critical and can be treated as a don't-care condition.

As a hint to guide your design process, consider utilizing the previously developed FSM tailored for the PS/2 packet parser and integrate a datapath capable of capturing and storing the incoming byte data. This combination will form the core functionality of the top_module you are tasked to implement. Keep in mind to design this module while adhering to a synchronous reset approach.