// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Given an 8-bit input vector [7:0], reverse its bit ordering.

//Hint: assign out[7:0] = in[0:7]; does not work because Verilog does not allow vector bit ordering to be flipped.
//The concatenation operator may save a bit of coding, allowing for 1 assign statement instead of 8.

module top_module( 
    input [7:0] in,
    output [7:0] out
);

	// Insert your code here
	
endmodule
