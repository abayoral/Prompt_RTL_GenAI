module top_module(
    input in,
    output out
);

    // Direct assignment to reflect wire behavior
    assign out = in;

endmodule