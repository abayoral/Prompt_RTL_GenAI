You hold the esteemed position of a senior Digital Design Engineer at a prestigious company specializing in advanced hardware design, and you have been entrusted with the formidable task of developing a crucial Verilog module for a cutting-edge product that is anticipated to be integral to your company's next-generation offerings. The success of this particular module is crucial not only for the innovative product's functionality but also for upholding and further enhancing your company's esteemed reputation within the highly competitive computer hardware industry.

The specific design requirement calls for the construction of a robust 32-bit global history shift register that is equipped with the capability to rollback its state when a pipeline flush is necessitated by a branch misprediction. This requires a precise mechanism capable of adjusting the history register dynamically.

In the scenario where a branch prediction is made, signaled by an active high signal `predict_valid` (i.e., `predict_valid = 1`), it is essential to update the branch history by shifting in the bit `predict_taken` at the least significant bit (LSB) side of the register. This shift effectively updates the branch history to reflect the predicted behavior, where `predict_history[0]` denotes the predicted direction of the most recently encountered (youngest) branch in terms of prediction.

Conversely, when a branch misprediction is detected, indicated by `train_mispredicted = 1`, it is crucial to reload the branch history register with the correct state as it should appear after completing the mispredicted branch. This involves loading a history that combines the preceding history prior to the misprediction (`train_history`) with the actual outcome of the branch (`train_taken`), which reflects the post-misprediction branch behavior accurately.

Notably, in situations where the signals for both a prediction and a misprediction are active concurrently, the misprediction must take priority. The rationale is that the pipeline flush initiated by the misprediction will also annul the effects of any current branch prediction that is simultaneously in process.

The `predict_history` output needs to effectively represent the current state of the branch history register. Additionally, there is an asynchronous reset signal, `areset`, that, when activated, must reset the entire history counter to zero, ensuring that the system returns to a consistent and known state.

Your task is to design and implement this module, named `top_module`, with the specified inputs and outputs that adhere to the described functionality and handle the aforementioned conditions efficiently. This entails dealing with edge cases correctly and ensuring that the module performs reliably under different operational states. Consider aspects such as timing, resource usage, and any potential hazards that might arise during its integration into the wider system.