As a senior Digital Logic Design Engineer at a prominent hardware design company, your responsibilities include the development of essential components for cutting-edge products. One of the most critical tasks you are currently facing involves designing a Verilog module that performs a specific function—namely, a "population count" circuit. The purpose of this circuit is to accurately tally the number of '1' bits present within a given input vector. This module is particularly significant as its successful implementation will play a key role in upholding the company's reputation within the competitive landscape of computer hardware design.

The requirement for this task involves creating a population count circuit tailored for a 3-bit input vector, which means the design must effectively process an input consisting of three bits and produce an output that accurately reflects the total count of '1's seen in that input. The output must be a 2-bit vector, as there can be a maximum of three '1' bits in a 3-bit input, which can be represented in binary form using 2 bits.

With that context in mind, the question is how to approach the design and implementation of this Verilog module. What considerations should be taken into account when developing a circuit that can reliably perform the population count for a 3-bit input vector? What design strategies, coding practices, and testing methodologies would ensure that the module functions correctly and meets the expectations for performance and reliability within your company's product?