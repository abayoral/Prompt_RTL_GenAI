
To build a comprehensive knowledge base for generating Verilog modules, consider the following categories of information: Verilog fundamentals, design principles, common patterns, debugging tips, and best practices. Here’s a detailed look into each category:

### Verilog Fundamentals
1. **Data Types**:
   - **Reg and Wire**: Understand the differences and appropriate use cases for `reg` and `wire`.
   - **Vectors**: Use vectors for groupings of bits (e.g., `[7:0]` for 8-bit wide data).
   - **Parameter**: Utilize parameters for defining constants and making modules configurable.

2. **Operators**:
   - **Logical vs. Bitwise**: Use logical operators (`&&`, `||`, `!`) for conditions and bitwise operators (`&`, `|`, `~`) for bit manipulation.
   - **Arithmetic**: Common arithmetic operators include `+` (addition), `-` (subtraction), `*` (multiplication), and `/` (division).

3. **Control Structures**:
   - **Always Blocks**: Difference between `always @(posedge clk)`, `always @(negedge clk)`, `always @*`, and others.
   - **Case Statements**: Proper usage and default cases for coverage.

4. **Modules and Hierarchy**: 
   - **Module Declaration**: Syntax for defining modules, inputs, outputs, and instantiating sub-modules.
   - **Hierarchy**: Understanding how modules interact and can be connected.

### Design Principles
1. **Synchronous vs. Asynchronous Design**:
   - **Clocked Logic**: Use synchronous design principles where state changes on clock edges.
   - **Reset Handling**: Incorporate asynchronous and synchronous resets in designs.

2. **Combinational vs. Sequential Logic**:
   - **Combinational Logic**: Designed using `always @*` without clocks.
   - **Sequential Logic**: Use `always @(posedge clk)` for stateful elements.

3. **Design for Synthesis (DFS)**:
   - Writing synthesizable code: Avoid system tasks/functions and ensure the logic is realizable in hardware.
   - **RTL Design**: Ensure proper register transfer level (RTL) coding styles that are synthesizable.

### Common Patterns
1. **State Machines**:
   - One-hot and binary encoding for state machines.
   - Encoding states properly and using `enum` for readability.

2. **Pipelining**: 
   - Techniques for pipeline stages to boost design performance.
   - Balancing register and combinational logic delays.

3. **Timing Constraints**:
   - Setup and hold time considerations.
   - Clock domain crossing (CDC) techniques to avoid metastability.

### Debugging Tips
1. **Simulation**:
   - Using testbenches, initial blocks, and display tasks for verifying functionality.
   - Understanding waveforms and timing diagrams for debugging.

2. **Linting and Formal Verification**:
   - Using linting tools to catch common mistakes and coding style violations.
   - Formal verification for checking properties and assertions.

3. **Common Bugs**:
   - Avoiding race conditions in combinational and sequential logic.
   - Proper signal initialization and reset.

### Best Practices
1. **Modular Design**:
   - Breaking down complex designs into smaller sub-modules.
   - Encapsulation, reusability, and maintainability of modules.

2. **Code Readability**:
   - Clear and consistent naming conventions for signals and modules.
   - Adequate commenting to clarify purpose and functionality of the code.

3. **Test Coverage**: 
   - Writing exhaustive testbenches to cover all possible scenarios.
   - Using random testing and corner cases to ensure robustness.

By comprehensively understanding these topics, a language model will be better equipped to generate efficient, reliable, and accurate Verilog modules for various digital design problems.

Task:
The following adder-subtractor with zero flag doesn't work. Fix the bug(s).


// synthesis verilog_input_version verilog_2001
module top_module ( 
    input do_sub,
    input [7:0] a,
    input [7:0] b,
    output reg [7:0] out,
    output reg result_is_zero
);//

    always @(*) begin
        case (do_sub)
          0: out = a+b;
          1: out = a-b;
        endcase

        if (~out)
            result_is_zero = 1;
    end

endmodule