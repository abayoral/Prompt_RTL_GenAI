module top_module(
    output one
);

// Assign a constant logic high value to the output signal
    assign one = 1'b1;

endmodule