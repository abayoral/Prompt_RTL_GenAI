// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Make a decade counter that counts 1 through 10, inclusive. The reset input is synchronous, and should reset the counter to 1.

module top_module (
    input clk,
    input reset,
    output [3:0] q);

    // Insert your code here

endmodule