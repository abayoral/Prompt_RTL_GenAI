// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Build a combinational circuit with 100 inputs, in[99:0].

// There are 3 outputs:

// out_and: output of a 100-input AND gate.
// out_or: output of a 100-input OR gate.
// out_xor: output of a 100-input XOR gate.

// Hint: The reduction operators will be useful here.

module top_module( 
    input [99:0] in,
    output out_and,
    output out_or,
    output out_xor 
);

	// Insert your code here

endmodule