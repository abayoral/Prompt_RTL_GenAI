module top_module( output one );

    // Assign constant logic high (1) to the output
    assign one = 1'b1;

endmodule