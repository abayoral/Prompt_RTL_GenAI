module top_module (
    output wire one
);
    // Assign logic high (1) to the output
    assign one = 1'b1;  // Using 1'b1 to explicitly denote 1 in binary format

endmodule