
### Verilog Design Background Knowledge

#### Verilog Language Basics
1. **Module Definition**: A Verilog module defines a hardware block. It consists of:
   - **Port Declaration**: Describes input and output signals.
   - **Internal Register/Wire Declaration**: Variables used within the module.
   - **Behavioral/Structural Code**: Describes what the module does, either behaviorally (using statements) or structurally (using other module instantiations).

2. **Data Types**
   - `reg`: Variable used to hold values in procedural blocks like `always`.
   - `wire`: Variable representing physical wires, used for continuous assignment or connections between modules.
   
3. **Procedural Blocks**:
   - **always block**: Executes whenever a specified event occurs, such as a change in clock or reset.
     - `always @ (posedge clk)`: Trigger on the positive edge of the clock.
     - `always @ (*)`: Trigger whenever any variable in the sensitivity list changes.

4. **Blocking vs Non-Blocking Assignments**:
   - `=`: Blocking assignment, used in combinational logic.
   - `<=`: Non-blocking assignment, used in sequential logic to ensure proper timing of updates.

#### Sequential Logic Design Principles
1. **Clocking and Timing**
   - Synchronous designs rely on clock signals to synchronize changes in state.
   - Asynchronous signals, such as reset, are not synchronized to the clock. Care must be taken to avoid metastability.

2. **Reset Logic**
   - **Asynchronous Reset**: Can reset the state of the module upon activation, independent of the clock.
   - **Synchronous Reset**: Resets the state in synchronization with the clock edge.

3. **Control Signals**
   - Enable signals (`ena`): Used to control whether certain operations occur, such as shifting in a shift register.
   - Load signals (`load`): Used to load specific data into the registers.

4. **Priority in Control Signals**
   - When multiple control signals are active simultaneously, priority must be defined to avoid conflicts. Typically, loading data has a higher priority than enabling another operation like shifting.

#### Common Constructs and Best Practices
1. **Shift Registers**
   - Sequential elements that shift their content left or right with each clock cycle.
   - Can include additional logic to load new data or reset the contents.

2. **Synchronous Load**
   - Loading data on the same clock edge can be prioritized by checking the load signal first, before any shifting or other operations.

3. **Verilog Code Structuring**
   - Use clear and descriptive signal names.
   - Encapsulate related logic in understandable blocks.
   - Maintain consistent formatting for readability and maintainability.

4. **Defensive Coding**
   - Always specify the full width of vectors.
   - Ensure sensitivity lists in always blocks are complete.
   - Careful handling of edge conditions and race conditions, especially with asynchronous resets.

### Principles for Verilog Design Enhancements

1. **Modularity and Reusability**
   - Design modules to be as modular and reusable as possible.
   - Keep functionalities well-encapsulated; avoid interdependencies that can make the module hard to reuse.

2. **Hierarchy and Abstraction**
   - Use hierarchical design to break complex designs into simpler, smaller modules.
   - Abstract details within lower-level modules, exposing upper levels only to necessary interfaces.

3. **Simulation and Testing**
   - Design with verification in mind. Write testbenches to validate functionalities before synthesizing hardware.
   - Use assertions to check for invariances and unexpected conditions during simulation.

4. **Resource Efficiency**
   - Implement designs that are resource-efficient. Optimize for area, power, and performance.
   - Use design constructs that appropriately map to the target technology (FPGA/ASIC).

5. **Documentation and Comments**
   - Thoroughly document functionality, inputs, outputs, and the role of each significant piece of logic.
   - Use comments to explain complex logic or unusual cases.

### Common Patterns in Verilog Design
1. **Finite State Machines (FSMs)**
   - Often used for control logic with clearly defined states and transitions.

2. **Pipelining**
   - Technique to achieve higher throughput by breaking operations into multiple clock-cycle stages.

3. **Clock Domain Crossing (CDC)**
   - Special care when transferring signals between different clock domains to avoid metastability.

4. **Parameterized Designs**
   - Use parameters to create flexible and scalable modules that can be easily configured.

### Summary
By understanding and applying these principles, knowledge, and best practices, language models can more effectively generate efficient, accurate, and maintainable Verilog code. This provides a comprehensive foundation that can enhance Verilog design tasks across a broad range of applications.

Task:
// Build a 4-bit shift register (right shift), with asynchronous reset, synchronous load, and enable.

// areset: Resets shift register to zero.
// load: Loads shift register with data[3:0] instead of shifting.
// ena: Shift right (q[3] becomes zero, q[0] is shifted out and disappears).
// q: The contents of the shift register.
// If both the load and ena inputs are asserted (1), the load input has higher priority.

module top_module(
    input clk,
    input areset,  // async active-high reset to zero
    input load,
    input ena,
    input [3:0] data,
    output reg [3:0] q); 


    // Insert your code here

endmodule
