Assume you are a seasoned Digital Design Engineer working at a highly respected hardware design firm. You have been assigned the critical task of creating a Verilog module that will play an essential role in the development of an advanced, next-generation product. The success of this particular module is vital for upholding the esteemed reputation of your company within the competitive computer hardware industry. 

Imagine you are working on the design of a digital circuit responsible for managing the ringer and vibration motor of a cell phone. When an incoming call is detected (indicated by the input signal `ring`), your circuit needs to decide between activating the phone's ringer (setting the output `ringer` to logical 1) or turning on the vibration motor (setting the output `motor` to logical 1), but importantly, it should not enable both simultaneously. 

If the phone is set to vibrate mode, as indicated by the input signal `vibrate_mode` being set to 1, your circuit should enable the vibration motor instead of the ringer. Conversely, if the vibrate mode is not active, the ringer should be activated.

The challenge is to implement this logic using Verilog, particularly focusing on utilizing assign statements. This involves translating the given problem description into a network of logic gates, ensuring the logic is accurately represented in hardware language. 

Consider approaching this problem with a mindset often used in hardware design which focuses on the desired state of outputs first and then traces back to the inputs that cause these states. Unlike traditional sequential programming approaches where the sequence of events is thought of as "If (inputs are ___), then (outputs should be ___)", in hardware design, the mindset shifts towards "The (output should be ___) when (inputs are ___)", starting from the desired condition of outputs and reasoning back to the necessary conditions of inputs.

In this scenario, reframe your logic thinking by considering conditions such as "The motor is active under the condition that ___" instead of framing it sequentially with "If the phone is in vibrate mode, then ___". 

In summary, translate this logic into a Verilog module using the assign statement methodology, ensuring that only one output is active at any time based on the input conditions, reflecting the operational needs of a phone's ringer and vibration system. Your task is to structure and implement this logic efficiently within the constraints of hardware design principles.