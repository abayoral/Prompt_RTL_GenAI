As a senior Digital Design Engineer at your company, you have been entrusted with the vital task of developing a Verilog module that serves as a gshare branch predictor for a cutting-edge hardware product. This module's performance and reliability are crucial for your organization's standing in the competitive computer hardware industry. Your objective is to construct a gshare branch predictor that operates based on a 7-bit program counter (PC) and a 7-bit global history register, which undergo a bitwise XOR operation to generate a 7-bit index. This index is then utilized to retrieve data from a pattern history table (PHT) composed of 128 two-bit saturating counters. The structure encompasses a 7-bit global branch history register.

The branch predictor operates with two distinct sets of interfaces. One interface handles the prediction process, utilized during the Fetch stage of the processor to provide branch direction forecasts for instructions being retrieved. The other interface is responsible for training, updating the predictor's accuracy based on determined branch outcomes as branch instructions are executed throughout the pipeline.

When a branch prediction is invoked (signaled by `predict_valid = 1`) for a specific program counter, the predictor must deliver both the anticipated branch direction and the current state of the branch history register utilized for the prediction. Upon the next positive clock edge, the branch history register is updated in response to the forecasted branch.

Conversely, when a training request is made (indicated by `train_valid = 1`), the predictor receives the program counter, the branch history register's value associated with the branch in question, the actual outcome of the branch, and whether there was a misprediction that necessitated a pipeline flush. The objective here is to adjust the PHT to enhance the predictor’s accuracy for similar branches in the future. Further, should the branch have been mispredicted, the predictor must also restore the branch history register to its configuration right after the errant branch's execution concluded.

In scenarios where both a training operation for a misprediction and a prediction request for a different, younger instruction occur simultaneously, the training is prioritized as the impending prediction will be rendered moot. When training and predicting the same PHT entry occur concurrently, the prediction accesses the initial PHT state predating the training, since adjustments to the PHT occur at the subsequent positive clock edge. An outlined timing diagram visually portrays how the system manages concurrent training and predictions on PHT entry 0 across cycles, illustrating that a training request in cycle 4 impacts the PHT only by cycle 5, while a simultaneous prediction request in cycle 4 remains unaffected by these changes.

Additionally, the system incorporates an asynchronous reset, denoted as `areset`, which uniformly resets the PHT to a default state of `2'b01` (interpreted as weakly not-taken) while clearing the global history register to zero.

Your goal is to integrate this design logic efficiently within the Verilog module, delineated as `top_module`, complete with its respective inputs and outputs. Through this, ensure comprehensive functionality so the branch predictor can accurately provide and adjust branch direction predictions, leveraging both the program counter and branch history register inputs for its operations.