As a Senior Digital Design Engineer at a leading hardware design company, you are assigned the crucial task of creating a Verilog module that functions as a gshare branch predictor for an upcoming next-generation product. The successful development of this module is of utmost importance, as it plays a vital role in sustaining your company's esteemed reputation within the competitive landscape of computer hardware design.

The primary goal of this task is to design a branch predictor that utilizes a 7-bit program counter (PC) alongside a 7-bit global history. This configuration will be hashed through an XOR operation to generate a 7-bit index, which will subsequently access a table consisting of 128 entries that each contain two-bit saturating counters. Additionally, the branch predictor must incorporate a global branch history register that is also 7 bits in size.

The branch predictor must facilitate two distinct sets of interfaces: one dedicated to making predictions and the other aimed at training the predictor itself. The prediction interface will be engaged during the processor's fetch stage, wherein it will request predictions regarding the direction of branches for the instructions currently being fetched. Following the execution of these branches, the actual outcomes will become available, allowing for the training of the branch predictor based on this real-time data. 

When a branch prediction is sought (indicated by `predict_valid` being set to 1) for a specified PC, the predictor should return both the predicted branch direction and the state of the branch history register utilized for this prediction. It is essential that the branch history register is updated at the next positive clock edge in accordance with the predicted branch.

In contrast, when a training request is made (indicated by `train_valid` being set to 1), the predictor needs to receive the current PC and the value of the branch history register related to the branch being trained, along with the actual outcome of the branch and a signal indicating whether there was a misprediction that necessitates a pipeline flush. The update process must include refining the pattern history table (PHT) to enhance the accuracy of future predictions for this particular branch. Moreover, if the training involves a misprediction, it is crucial to restore the branch history register to the state it was in immediately following the execution of the mispredicted branch.

A complex situation arises when both prediction and training requests occur in the same cycle. In such cases, priority is given to the training operation, as the predicted branch is ultimately irrelevant if it involves a misprediction. If both prediction and training of the same PHT entry happen simultaneously, it is important to recognize that the prediction sees the state of the PHT before the training takes effect, which happens only on the next positive clock edge.

Lastly, it’s worth noting that an asynchronous reset (`areset`) is incorporated into the design, serving to clear the entire PHT to a default state of 2b'01 (weakly not-taken) and resetting the global history register to zero.

With this understanding, the question at hand is: How can you effectively implement this gshare branch predictor in Verilog, ensuring that all specified functionalities, timing considerations, and operational priorities are properly addressed within the module structure provided?