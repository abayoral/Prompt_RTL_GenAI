// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Create a 100-bit binary adder. The adder adds two 100-bit numbers and a carry-in to produce a 100-bit sum and carry out.

// Hint: There are too many full adders to instantiate, but behavioural code works in this case.

module top_module( 
    input [99:0] a, b,
    input cin,
    output cout,
    output [99:0] sum );

    // Insert your code here

endmodule

