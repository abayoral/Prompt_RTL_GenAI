module top_module (
    input wire in,   // Input signal
    output wire out  // Output signal
);
    // Direct wire connection
    assign out = in;
endmodule