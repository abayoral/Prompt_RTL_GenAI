// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Create a module that implements a NOR gate. 
// A NOR gate is an OR gate with its output inverted. 
// A NOR function needs two operators when written in Verilog.

// Hint: Verilog has separate bitwise-OR (|) and logical-OR (||) operators, like C. 
// Since we're working with a one-bit here, it doesn't matter which we choose.

module top_module( 
    input a, 
    input b, 
    output out );

// Insert your code here

endmodule
