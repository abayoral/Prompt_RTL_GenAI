// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Create a module that implements a NOT gate.

//Hint: Verilog has separate bitwise-NOT (~) and logical-NOT (!) operators, 
//like C. Since we're working with a one-bit here, it doesn't matter which we choose.

module top_module( input in, output out );

//Insert your code here

endmodule
