
### Verilog Design Knowledgebase

#### General Concepts

1. **Hierarchical Design**:
   - Break down complex designs into smaller, manageable modules.
   - Use hierarchical design to encapsulate functionality and promote reuse.

2. **Data Types**:
   - **Wire**: Used to connect different components and represent combinational logic.
   - **Reg**: Used to store values and represent sequential logic.
   - **Vector**: Multiple-bit wires or registers (e.g., `[15:0]`).

3. **Structural vs. Behavioral Modeling**:
   - **Structural**: Using instantiation of modules to build a design.
   - **Behavioral**: Using high-level constructs (e.g., `always` blocks, `case` statements).

4. **Sensitivity List**:
   - Defines when a block of code should be evaluated.
   - Commonly uses `always @(*)` for combinational logic and `always @(posedge clk)` for sequential logic.

5. **Blocking and Non-Blocking Assignments**:
   - **Blocking (`=`)**: Executes statements sequentially within an `always` block.
   - **Non-Blocking (`<=`)**: Allows statements to execute concurrently, typically used in sequential logic.

#### Principles and Best Practices

1. **Modular Design**:
   - Encapsulate functionality within modules.
   - Interface modules using well-defined `input` and `output` ports.

2. **Coding Style Guidelines**:
   - Use meaningful names for ports and signals.
   - Comment code sufficiently for readability and maintenance.
   - Maintain consistent indentation and formatting.

3. **Synchronization**:
   - Handle asynchronous inputs carefully to avoid metastability.
   - Use synchronization registers for clock domain crossing.

4. **State Machines**:
   - Design state machines with clear state encoding.
   - Use `case` statements for readability and maintainability.
   - Define default states to handle unexpected conditions.

5. **Testbenches**:
   - Develop comprehensive testbenches to validate functionality.
   - Include test cases for normal, boundary, and exceptional conditions.
   - Use assertions where applicable for automatic checking of conditions.

#### Common Patterns

1. **Mux (Multiplexer)**:
   - Use a `case` statement to switch between different inputs based on a selector.
   - Example: A 9-to-1 mux selecting between nine 16-bit inputs.

2. **Decoder**:
   - Decode binary inputs into a one-hot representation.
   - Common for address decoding and selecting specific lines.

3. **Encoders**:
   - Encode multiple input lines into a smaller binary representation.
   - Often used in priority encoding and interrupt handling.

4. **Flip-Flops and Latches**:
   - Use `always @(posedge clk)` for flip-flops.
   - Use `always @(*)` or `if` statements for latches, but avoid due to potential unintended latches.

5. **Finite State Machines (FSMs)**:
   - Define states and transitions clearly.
   - Use `parameter` to define state values for clarity.

#### Example Principles for Mux Implementation

1. **Case Statement Usage**:
   - A `case` statement is ideal for selecting between multiple inputs based on a selector value.
   - Ensure all cases are covered, and provide a default case for unexpected values.

2. **Default Output**:
   - For unused selector values, define a default output (e.g., all `1`s for `sel` values 9 to 15).

3. **Parameterization**:
   - Consider using parameters to make the design scalable and reusable.

### Applying These Principles

- **Selector Range**: Include 9 to 15 in the `case` statement to handle default values.
- **Combinational Logic**: Use `always @(*)` for combinational selection logic.
- **Output Initialization**: Ensure the output is initialized, especially for default cases.
- **Comments and Clarity**: Maintain clear, expressive comments throughout the code for maintainability.

By utilizing these principles and common patterns, Verilog design tasks such as creating a multiplexer can be executed effectively, ensuring robust and maintainable code.

Task:
// Create a 16-bit wide, 9-to-1 multiplexer. sel=0 chooses a, sel=1 chooses b, etc. 
// For the unused cases (sel=9 to 15), set all output bits to '1'.

// Hint: With this many options, a case statement may be useful.

module top_module( 
    input [15:0] a, b, c, d, e, f, g, h, i,
    input [3:0] sel,
    output [15:0] out );

    //Insert your code here

endmodule