In your role as a senior Digital Design Engineer at a prominent hardware design company, you have been entrusted with the development of an essential Verilog module that plays a crucial role in the rollout of a next-generation product. The company’s reputation within the competitive computer hardware industry hinges on the success of this module, making its design and operation vital.

Your task is to design a priority encoder for 8-bit inputs. The objective of this module is to intake an 8-bit vector and successfully identify and report the index of the first '1' bit starting from the least significant bit position. If the vector contains no bits set to '1', the output should return zero. It is imperative to ensure that the design meets this functionality accurately, as incorrect reporting of bits could have significant repercussions on the product's performance.

For example, consider the input vector 8'b10010000. In this scenario, the priority encoder should output the decimal value 4, expressed as a 3-bit binary 3'd4, because the first '1' encountered from the right-hand side (starting from bit[0]) is at position bit[4].

Additionally, you are required to adhere to the Verilog 2001 standard, which imposes specific syntax and design practices, ensuring compatibility and synthesis readiness across various tools that support this version of Verilog.