As a senior Digital Design Engineer actively involved in hardware development, you are faced with the task of designing a crucial Verilog module that is essential for an upcoming next-generation product. The successful implementation of this module is not just a technical requirement; it carries significant implications for upholding the reputation and competitiveness of your computer hardware company within the industry.

Your specific objective is to construct a finite-state machine (FSM) that is capable of detecting a predefined sequence, specifically the bit sequence '1101', within a continuous stream of input bits. Upon successful detection of this sequence, the FSM must set a particular output signal, `start_shifting`, to a high state (1), and maintain this state indefinitely until it receives a reset signal. It is important to note that the FSM is designed to remain in this final state purposefully; this design choice is intended to model the transition to additional states that will be incorporated into a more comprehensive FSM in subsequent development exercises.

With the design constraints and the intended functionality in mind, you are tasked with creating an appropriate module structure in Verilog. The module, referred to as `top_module`, includes inputs for a clock signal (`clk`), a synchronous reset signal (`reset`), and a data input signal (`data`). It also includes an output signal (`start_shifting`) that indicates the successful detection of the sequence. 

In light of this context, what specific considerations and strategies should be employed in the design of the FSM to ensure that it effectively and efficiently detects the sequence '1101'? Additionally, what best practices should be followed in the Verilog code implementation to facilitate future extensions of the FSM's capabilities as envisioned in the upcoming development phases?