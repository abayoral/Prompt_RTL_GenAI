// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Implement the following D flip-flop with asynchronous reset

module top_module (
    input clk,
    input d, 
    input ar,   // asynchronous reset
    output q);

    // Insert your code here

endmodule


