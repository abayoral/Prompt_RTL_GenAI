
### Verilog Knowledge Base for Language Model

#### Fundamental Concepts and Terminologies

1. **Modules and Ports:**
   - A module in Verilog is a fundamental building block.
   - Modules have input and output ports used for communication with other modules.
   - Ports are declared with `input`, `output`, or `inout`.

2. **Data Types:**
   - Basic data types: `wire`, `reg`, `integer`, `real`.
   - `wire` is used for combinational logic.
   - `reg` is used for storage elements like flip-flops.

3. **Operators:**
   - Arithmetic operators: `+`, `-`, `*`, `/`
   - Relational operators: `==`, `!=`, `<`, `>`, `<=`, `>=`
   - Logical operators: `&&`, `||`, `!`
   - Bitwise operators: `&`, `|`, `^`, `~`

4. **Gate-Level Modeling:**
   - Basic gates: `and`, `or`, `not`, `nand`, `nor`, `xor`, `xnor`.

5. **Combinational and Sequential Logic:**
   - **Combinational Logic:** Output depends only on the current inputs. Examples include adders, multiplexers, etc.
   - **Sequential Logic:** Output depends on the current inputs and the past history (state). Examples include flip-flops, counters, etc.

6. **Blocking vs Non-blocking Assignments:**
   - Blocking (`=`): Executes statements sequentially within initial or always blocks.
   - Non-blocking (`<=`): Executes statements concurrently within always blocks.

7. **Always Blocks:**
   - Used to describe both combinational and sequential logic.
   - `always @*`: Represents combinational logic.
   - `always @(posedge clk)` or `always @(negedge clk)`: Represents sequential logic triggered by clock edges.

8. **Sensitivity List:**
   - List of signals that trigger the execution of an `always` block.
   - `always @*` is a shorthand for "whenever any input changes".

#### Principles and Best Practices

1. **Consistent Naming Conventions:**
   - Use meaningful and consistent names for signals, modules, and variables.

2. **Structured Design:**
   - Break complex designs into smaller, reusable submodules.
   - Follow a hierarchical modeling approach to maintain clarity.

3. **Coding for Synthesis:**
   - Ensure the code can be synthesized into hardware respecting timing and resource constraints.
   - Avoid constructs that are not synthesizable (e.g., delays, real numbers).

4. **Testbenches:**
   - Develop testbenches to simulate and verify the functionality of your design.
   - Include all possible input scenarios, including edge cases.

5. **RTL Design Patterns:**

   - **Adder/Subtractor:**
     - Use simple constructs like `assign` for combinational adders.
     - Ensure correct management of carry bits.

   - **State Machines:**
     - Use `case` or `if-else` statements to model state transitions.
     - Use enumerations for state encoding.

   - **Decoders/Encoders:**
     - Use `always @*` to describe combinational logic of encoders and decoders.
   
   - **Multiplexers:**
     - Use `always @*` or `assign` to describe the selection logic.

6. **Common Practices for Full Adders:**
   - A full adder adds three binary bits (A, B, Cin) and produces a Sum and Cout.
   - The Cout is used as a carry-in for the next stage if chaining multiple adders.

7. **Modular Design:**
   - Always design with reusability in mind.
   - Modular designs help in easier debugging and testing.

### Common Patterns

1. **Adder Pattern:**
   - **Half Adder:** Produces sum and carry from two bits.
   - **Full Adder:** Extends half adder to include carry-in.

2. **Multiplexer Pattern:**
   - Selects one of several input signals based on select lines.

3. **Flip-Flop Pattern:**
   - Basic memory element that stores a single bit, triggered by clock edges.

4. **Counter Pattern:**
   - Sequential circuit that counts upwards or downwards based on clock and control inputs.

5. **State Machine Pattern:**
   - Describes the behavior of sequential logic systems that transition between different states.

### Documentation and Comments

1. **Inline Comments:**
   - Use `//` for single-line comments to explain logic and important lines.

2. **Block Comments:**
   - Use `/* ... */` for multiline comments providing detailed descriptions or sections of the code.

3. **Port Descriptions:**
   - Clearly describe the role of each port in terms of the system’s functionality.

### Example Theoretical Explanation

For a Full Adder:
- **Inputs:**
  - `a`: First bit input.
  - `b`: Second bit input.
  - `cin`: Carry input from previous stage.
- **Outputs:**
  - `sum`: Sum output of `a`, `b`, and `cin`.
  - `cout`: Carry output to the next higher-order bit.

Understanding these fundamental principles and concepts aids in adhering to best practices, improving modularity, reusability, and maintainability of Verilog designs.

Task:
//Create a full adder. A full adder adds three bits (including carry-in) and produces a sum and carry-out.

module top_module( 
    input a, b, cin,
    output cout, sum );

    // Insert your code here

endmodule
