// you're a senior FPGA Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Implement the following circuit:

// in --- out

module top_module (
    input in,
    output out);
    
    // Insert your code here
endmodule
