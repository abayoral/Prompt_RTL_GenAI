// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Create a module that implements an AND gate.

// Hint: Verilog has separate bitwise-AND (&) and logical-AND (&&) operators, like C. 
// Since we're working with a one-bit here, it doesn't matter which we choose.

module top_module( 
    input a, 
    input b, 
    output out );

// Insert your code here

endmodule
