// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

//Create a module that implements an XNOR gate.

//Hint: The bitwise-XOR operator is ^. There is no logical-XOR operator.

module top_module( 
    input a, 
    input b, 
    output out );

// Insert your code here

endmodule
