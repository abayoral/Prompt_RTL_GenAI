// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Create a circuit that has two 2-bit inputs A[1:0] and B[1:0], and produces an output z. 
// The value of z should be 1 if A = B, otherwise z should be 0.


module top_module ( input [1:0] A, input [1:0] B, output z ); 
	// Insert your code here
endmodule
