// you're a senior Logic Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining the company's reputation in the industry.

// The 7458 is a chip with four AND gates and two OR gates. 

// Create a module with the same functionality as the 7458 chip. 
// It has 10 inputs and 2 outputs. You may choose to use an assign statement 
// to drive each of the output wires, or you may choose to declare (four) wires 
// for use as intermediate signals, where each internal wire is driven by the 
// output of one of the AND gates. For extra practice, try it both ways.


// Hint: You need to drive two signals (p1y and p2y) with a value.

module top_module ( 
    input p1a, p1b, p1c, p1d, p1e, p1f,
    output p1y,
    input p2a, p2b, p2c, p2d,
    output p2y );

// Insert your code here

endmodule