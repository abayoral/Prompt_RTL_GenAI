module top_module(
    output wire zero
);
    // Assign the constant value 0 to the output zero
    assign zero = 1'b0;
endmodule