// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

//Build a circuit that has one 3-bit input, then outputs the same vector, 
// and also splits it into three separate 1-bit outputs. 
// Connect output o0 to the input vector's position 0, o1 to position 1, etc.

module top_module ( 
    input wire [2:0] vec,
    output wire [2:0] outv,
    output wire o2,
    output wire o1,
    output wire o0  ); // Module body starts after module declaration

// Insert your code here

endmodule
