// you're a senior hardware engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining the company's reputation in the industry.

//Build a combinational circuit with two inputs, a and b.

//There are 7 outputs, each with a logic gate driving it:

//out_and: a and b
//out_or: a or b
//out_xor: a xor b
//out_nand: a nand b
//out_nor: a nor b
//out_xnor: a xnor b
//out_anotb: a and-not b

module top_module( 
    input a, b,
    output out_and,
    output out_or,
    output out_xor,
    output out_nand,
    output out_nor,
    output out_xnor,
    output out_anotb
);
	// Insert your code here
endmodule
