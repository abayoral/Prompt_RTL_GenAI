We aim to enhance a serial receiver by incorporating a parity checking mechanism. In this context, parity checking involves appending an additional bit following each transmitted data byte. Specifically, we will employ odd parity, meaning the aggregate number of '1' bits across the total of 9 bits received (including the parity bit) should be odd. For instance, a sequence like `101001011` adheres to odd parity since it contains 5 '1' bits, whereas a sequence like `001001011` does not comply as it contains 4 '1' bits.

To achieve this, you are required to adapt both your finite state machine (FSM) and datapath to facilitate odd parity verification. The `done` signal should assert exclusively when a byte is correctly received, and it passes the parity check. The FSM should possess the capability, akin to the serial receiver FSM, to detect the start bit, monitor for all 9 bits comprising both the data and the parity, and then verify the correctness of the stop bit. Should the expected stop bit fail to appear in sequence, the FSM must seek out the subsequent occurrence of a stop bit before attempting to capture the next byte.

You have access to a module crafted for parity calculation from the input stream. This module, functioning as a Toggle Flip-Flop (TFF) equipped with a reset option, is designed to tally the number of '1' bits within each byte. It operates such that upon clocking, if reset is active, it sets the output `odd` to zero. Conversely, if the input is '1', it toggles the `odd` output.

Consider that the serial communication protocol proceeds by sending the least significant bit (LSB) initially, followed by the parity bit after the sequence of 8 data bits. Utilizing the given `parity` module, adapt your existing FSM and datapath architecture (from a baseline such as `Fsm_serialdata`) to incorporate the newly required functionality for parity checking in the `top_module`. Make sure to manage the sequence control and verification processes to affirm the integrity and correctness of each received byte after applying the parity check.