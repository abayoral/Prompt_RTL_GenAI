Imagine you are serving as a senior Digital Design Engineer at a prominent hardware design firm, and you have been assigned the important task of developing a critical Verilog module for a next-generation product. This module plays a key role in the overall functionality of the product and is crucial for preserving the company’s esteemed reputation within the competitive landscape of computer hardware design.

In this context, consider the design of a finite state machine (FSM) that is specifically intended to manage the operations of a motor. This FSM receives two types of inputs—labeled as x and y—originating from the motor, and it is responsible for producing two outputs, f and g, which directly influence the motor's operation. Additionally, the FSM is governed by a clock input, clk, and it features a reset input, resetn, which operates in an active-low manner.

The functional requirements of the FSM are as follows: while the reset input is asserted (active), the FSM must remain in an initial state, designated as state A. Once the reset signal is de-asserted, the FSM is expected to transition, after the next clock edge, and set the output f to 1 for a duration of one clock cycle. At this point, the FSM is required to begin monitoring the x input. Specifically, when x produces the sequence of values 1, 0, 1 over three consecutive clock cycles, the FSM should then transition to set the output g to 1 on the subsequent clock cycle.

While g remains at a value of 1, the FSM must continue to track the y input. If the y input registers a value of 1 within a maximum of two additional clock cycles, the FSM should ensure that g remains indefinitely at 1 (that is, it should persist in this state until a reset occurs). Conversely, if the y input does not receive a value of 1 within the stipulated two clock cycles, the FSM is to set g to 0 permanently (again, this state remains until reset).

Your challenge, therefore, is to implement this finite state machine correctly within the provided Verilog module structure. Taking into consideration the defined behavior and requirements, how would you approach the task of coding this FSM? What factors and design aspects would you prioritize in your implementation, and how would you ensure that all functional requirements are met? 

With the specifications laid out clearly, what design considerations will guide your development process, and what testing or validation methods will you employ to confirm that the FSM meets its operational criteria?