// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Module A is supposed to implement the function z = (x^y) & x. Implement this module.


module top_module (input x, input y, output z);

	// Insert your code here

endmodule
