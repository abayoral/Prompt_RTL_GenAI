module top_module( 
    input a, b, cin,
    output cout, sum );

    assign sum = a ^ b ^ cin; // Sum is XOR of a, b and cin
    assign cout = (a & b) | (b & cin) | (cin & a); // Carry out is when any two of the inputs are 1

endmodule