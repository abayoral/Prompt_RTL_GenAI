// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

//Build a circuit with no inputs and one output. That output should always drive 1 (or logic high).


module top_module( output one );

// Insert your code here
    assign one = [fixme];

endmodule
