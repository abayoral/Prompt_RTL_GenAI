// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Create 8 D flip-flops with active high asynchronous reset. All DFFs should be triggered by the positive edge of clk.

// Hint: The only difference in code between synchronous and asynchronous reset flip-flops is in the sensitivity list.

module top_module (
    input clk,
    input areset,   // active high asynchronous reset
    input [7:0] d,
    output [7:0] q
);

	// Insert your code here

endmodule
