
## Knowledge Base for Verilog Design

### Background Knowledge

1. **Introduction to Verilog:**
   - Verilog is a hardware description language (HDL) used to model electronic systems.
   - It allows designers to describe the behavior and structure of electronic circuits, especially digital logic circuits.

2. **Verilog Design Components:**
   - **Modules:** Basic building blocks in Verilog. They can represent anything from simple gates to complex processors.
   - **Ports:** Interfaces for modules. Ports are inputs and outputs through which a module communicates with the external world.
   - **Nets and Registers:** Nets represent connections between hardware elements (e.g., `wire`), while registers are variables that store values (e.g., `reg`).

### Principles of Verilog Design

1. **Hierarchical Design:** 
   - Break down complex systems into smaller, manageable modules.
   - Encourage modular design to improve readability and reusability.

2. **Parameterization:**
   - Use parameters to create reusable and configurable modules.
   - Parameters can define characteristics such as bit-widths, enabling modules to be adaptable for various applications.

3. **Clocking and Synchronization:**
   - Ensure proper synchronization in sequential circuits using clocks.
   - Consider clock domains and crossing when dealing with multiple clocks.

4. **Finite State Machines (FSM):**
   - Efficient way to model sequential logic.
   - Consists of states, transitions, and outputs based on current state and inputs.

5. **Testbenches:**
   - Crucial for verifying the functionality of your design.
   - Include stimulus generation, monitoring, and checking mechanisms.

### Best Practices

1. **Coding Conventions:**
   - Use clear and consistent naming conventions.
   - Comment your code to explain logic, especially complex sections.
   - Group related signals together (e.g., `input`, `output` declarations).

2. **Design for Testability:**
   - Include features that make it easy to test and debug.
   - Consider boundary cases and edge conditions in your design.

3. **Resource Optimization:**
   - Optimize for area, speed, and power depending on requirements.
   - Avoid unnecessary logic and redundant calculations.

4. **Use Behavioral Modeling:**
   - For complex combinational and sequential logic, behavioral modeling is often more succinct and easier to manage.
   - Behavioral modeling can be done using `always` blocks.

5. **Avoid Common Pitfalls:**
   - Ensure that all signals used in `always` blocks are appropriately declared as `reg`.
   - Avoid race conditions by writing deterministic code.
   - Ensure proper reset strategies for sequential circuits.

### Common Patterns in Verilog Design

1. **Adder/Subtractor:**
   - Describe using behavioral code to simplify the design.
   - Use conditional operator for handling carry and overflow in large bit-width scenarios.

2. **Registers and Flip-Flops:**
   - Utilize `always @(posedge clk)` for synchronous logic.
   - Handle asynchronous and synchronous resets correctly.

3. **Multiplexers:**
   - Use conditional operators (`? :`) or `case` statements for cleaner implementation.

4. **State Machines:**
   - Clearly define state encodings and transitions.
   - Use enumerated types (in SystemVerilog) for readability.

5. **Memory Elements:**
   - Leverage `reg [width-1:0]` arrays for memory representation.
   - Avoid combinational loops by ensuring memory reads occur in sequential logic blocks.

By incorporating these foundational concepts, principles, and patterns, another language model should have a robust knowledge base to generate high-quality Verilog modules suitable for various applications.

Task:
// Create a 100-bit binary adder. The adder adds two 100-bit numbers and a carry-in to produce a 100-bit sum and carry out.

// Hint: There are too many full adders to instantiate, but behavioural code works in this case.

module top_module( 
    input [99:0] a, b,
    input cin,
    output cout,
    output [99:0] sum );

    // Insert your code here

endmodule

