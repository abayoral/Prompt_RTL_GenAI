Imagine you are a seasoned Digital Design Engineer at a prominent hardware design company. Your responsibility is to develop a critical Verilog module that will serve as a key component in a next-generation product. The overall success and reputation of your company depend on the flawless implementation of this module.

Your task is to design a one-bit wide, 2-to-1 multiplexer. The multiplexer should operate such that when the select signal (sel) is 0, it outputs the value of input a; when sel is 1, it outputs the value of input b.

Consider using the ternary operator (formatted as condition ? value_if_true : value_if_false) to simplify your implementation and enhance code readability.

Below is the module outline provided as a starting point:

-----------------------------------------------------
module top_module( 
    input a, b, sel,
    output out 
); 

    // Insert your Verilog code implementation here

endmodule
-----------------------------------------------------

Your rephrased challenge is to create and complete the Verilog code for this multiplexer according to the specifications detailed above, ensuring that the routing of the input signals based on the select signal is correctly implemented. Keep the focus on clarity, readability, and adherence to the functional requirements as described.