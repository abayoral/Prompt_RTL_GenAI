// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Create 8 D flip-flops. All DFFs should be triggered by the positive edge of clk.

module top_module (
    input clk,
    input [7:0] d,
    output [7:0] q
);
	// Insert your code here

endmodule
