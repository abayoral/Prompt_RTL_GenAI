// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Build a 4-bit priority encoder. For this problem, if none of the input bits are high 
// (i.e., input is zero), output zero. Note that a 4-bit number has 16 possible combinations.

// Hint: Using hexadecimal (4'hb) or decimal (4'd11) number literals would save typing vs. binary (4'b1011) literals.

// synthesis verilog_input_version verilog_2001
module top_module (
    input [3:0] in,
    output reg [1:0] pos  );

    // Insert your code here

endmodule

