// you're a senior Digital Logic Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

//Build a circuit with no inputs and one output that outputs a constant 0
module top_module(
    output zero
);// Module body starts after semicolon

endmodule
