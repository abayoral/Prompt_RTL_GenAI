
## Knowledgebase for Verilog Design Tasks

### Fundamental Concepts
1. **Hardware Description Languages (HDLs)**: Understand that Verilog is an HDL used for describing electronic circuits and systems.

2. **Modules**: The primary building blocks in Verilog, similar to functions or classes in other programming languages. A module has an interface (with ports) and an internal structure.

3. **Port Declaration**: Ports define the inputs and outputs of a module. Generally, inputs, outputs, and inouts are declared at the top of the module.

4. **Registers and Wires**:
   - **reg**: Used for variables that hold values.
   - **wire**: Used for connecting different components.
   - **logic**: Preferred in SystemVerilog as it can act as both reg and wire.

5. **Always Blocks**: Used to describe behavior that changes over time, either synchronously (`always @(posedge clk)`) or asynchronously (`always @*`).

6. **Initial Blocks**: Used for initialization in simulation models.

7. **Assign Statements**: Continuous assignments used outside always blocks for combinational logic.

8. **Parameters**: Constants that can be defined for use within modules, making designs more customizable.

### Best Practices
1. **Modular Design**: Break down complex designs into smaller sub-modules for better readability and reusability.

2. **Naming Conventions**: Use clear and consistent naming for signals and modules to enhance readability and maintenance.

3. **Use of Comments**: Comment your code to explain non-obvious parts, particularly to clarify the intent of complex logic.

4. **Parameterized Designs**: Use parameters to create more flexible and reusable modules.

5. **Simulation and Testing**: Regularly simulate and test your design with different test cases to verify functionality.

### Common Patterns in Verilog Design
1. **Synchronous Logic**: Use `always @(posedge clk)` for describing logic that updates on clock edges.

2. **Asynchronous Reset**: Implementing reset functionality that initializes or resets the state of the system.
   ```verilog
   always @(posedge clk or posedge reset) begin
       if (reset) begin
           // reset logic
       end else begin
           // normal operation logic
       end
   end
   ```

3. **Finite State Machines (FSMs)**: Often used to control the sequential behavior of systems.
   - **State Encoding**: Use `enum` for state definitions in SystemVerilog.
   - **State Transition**: Next state logic and output logic within always blocks.

4. **Data Storage and Movement**: Use arrays and registers for storing and manipulating data.

5. **Bitwise Operations**: Efficiently use bitwise operations (`&`, `|`, `^`, `~`) for manipulating bits in registers and wires.

### Specific Concepts for Conway's Game of Life Implementation

1. **Grid Representation**: Think of the grid as a 2D array. In Verilog, this can be represented with a 1D array for simplicity:
   - A 16x16 grid can be represented as a `256-bit` vector.

2. **Neighbor Calculation**: For each cell, compute the number of live neighbors. This involves accessing the surrounding cells in the array:
   - Use modular arithmetic to handle the toroidal (wrap-around) property.

3. **State Transition Logic**: Given the rules of the game, implement the logic that transitions the state from one step to the next.

4. **Clock-Based Updates**: Ensure the system updates the grid state on each clock cycle:
   ```verilog
   always @(posedge clk) begin
       if (load) begin
           // load initial data into grid
       end else begin
           // update grid based on rules
       end
   end
   ```

5. **Loading Initial State**: Implement loading functionality to initialize the grid state from an external source or input vector.

### Additional Tools and Techniques
1. **Simulation Tools**: Use simulation tools like ModelSim or Vivado for testing and verifying your design.

2. **Synthesis Considerations**: Ensure that the design is synthesizable if the end goal is hardware implementation.

3. **Optimization**: Optimize logic for area, speed, and power consumption if designing for constrained environments.

4. **Version Control**: Use version control systems like Git for managing changes and collaboration on large projects.

By incorporating these principles, patterns, and best practices, a language model can generate more robust, efficient, and maintainable Verilog modules.

Task:
// Conway's Game of Life is a two-dimensional cellular automaton.

// The "game" is played on a two-dimensional grid of cells, where each cell is either 1 (alive) or 0 (dead). At each time step, each cell changes state depending on how many neighbours it has:

// 0-1 neighbour: Cell becomes 0.
// 2 neighbours: Cell state does not change.
// 3 neighbours: Cell becomes 1.
// 4+ neighbours: Cell becomes 0.
// The game is formulated for an infinite grid. In this circuit, we will use a 16x16 grid. To make things more interesting, we will use a 16x16 toroid, where the sides wrap around to the other side of the grid. For example, the corner cell (0,0) has 8 neighbours: (15,1), (15,0), (15,15), (0,1), (0,15), (1,1), (1,0), and (1,15). The 16x16 grid is represented by a length 256 vector, where each row of 16 cells is represented by a sub-vector: q[15:0] is row 0, q[31:16] is row 1, etc. (This tool accepts SystemVerilog, so you may use 2D vectors if you wish.)

// load: Loads data into q at the next clock edge, for loading initial state.
// q: The 16x16 current state of the game, updated every clock cycle.
// The game state should advance by one timestep every clock cycle.

// Hint: A test case that's easily understandable and tests some boundary conditions is the blinker 256'h7. It is 3 cells in row 0 columns 0-2. It oscillates between a row of 3 cells and a column of 3 cells (in column 1, rows 15, 0, and 1).

module top_module(
    input clk,
    input load,
    input [255:0] data,
    output [255:0] q ); 

    // Insert your code here

endmodule