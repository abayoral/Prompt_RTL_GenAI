module top_module(
    input a,
    input b,
    input c,
    output out
); 

    // Simplified expression from the Karnaugh map: the output is always 1
    assign out = 1;

endmodule