// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Build a circuit that will reverse the byte ordering of the 4-byte word.

// Hint: Part-select can be used on both the left side and right side of an assignment.
// AaaaaaaaBbbbbbbbCcccccccDddddddd => DdddddddCcccccccBbbbbbbbAaaaaaaa

module top_module( 
    input [31:0] in,
    output [31:0] out );

    //Insert your code here
    // assign out[31:24] = ...;

endmodule