// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

//Create a one-bit wide, 2-to-1 multiplexer. When sel=0, choose a. When sel=1, choose b.

//Hint: The ternary operator (cond ? iftrue : iffalse) is easier to read.

module top_module( 
    input a, b, sel,
    output out ); 

    // Insert your code here

endmodule
