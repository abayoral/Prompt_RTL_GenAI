module top_module(
    output wire one
);
    // Assign logic high (1) to the output
    assign one = 1'b1;
endmodule