module top_module ( 
    input p1a, p1b, p1c, p1d, p1e, p1f,
    output p1y,
    input p2a, p2b, p2c, p2d,
    output p2y );

    // Intermediate wires for AND gate outputs
    wire and1_out, and2_out, and3_out, and4_out;

    // AND gates for p1y
    assign and1_out = p1a & p1b & p1c; // First AND gate for p1y
    assign and2_out = p1d & p1e & p1f; // Second AND gate for p1y

    // AND gates for p2y
    assign and3_out = p2a & p2b; // First AND gate for p2y
    assign and4_out = p2c & p2d; // Second AND gate for p2y

    // OR gates for final outputs
    assign p1y = and1_out | and2_out; // OR gate for p1y
    assign p2y = and3_out | and4_out; // OR gate for p2y

endmodule