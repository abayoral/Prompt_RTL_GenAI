
### Verilog Design Knowledge Base

#### 1. **Verilog Fundamentals**
1. **Modules**:
   - The basic building blocks of Verilog designs. Encapsulate functionality and abstraction of digital circuits.
   - Defined using `module` and `endmodule` keywords.
   - Contains inputs, outputs, internal signals, and design logic.

2. **Data Types**:
   - **Nets (`wire`)**: Represent connections between hardware elements. Default data type used for passive signal propagation.
   - **Registers (`reg`)**: Used for variables that hold values between assignments, typically in procedural blocks (`always`, `initial`).

3. **Operators and Literals**: 
   - **Bitwise Operators**: `&` (AND), `|` (OR), `^` (XOR), `~` (NOT).
   - **Logical Operators**: `&&` (AND), `||` (OR), `!` (NOT).
   - **Number Literals**: Can be specified in binary (`4'b1010`), octal (`3'o7`), decimal (`4'd10`), or hexadecimal (`4'hA`).

#### 2. **Combinational Logic Design**
1. **Continuous Assignment**:
   - Using the `assign` keyword, continuously evaluates and assigns values to `wire` types.
   - Syntax: `assign <wire> = <expression>;`.

2. **Procedural Blocks**:
   - `always` blocks are used to describe both sequential and combinational logic.
   - `sensitive list` (`@`): Determines when the block executes.
     - Example for combinational logic: `always @(*)`.

3. **Priority Logic**:
   - Priority logic selects signals based on a hierarchy or precedence.
   - Can be implemented using `if-else` or `case` statements inside `always` blocks.

#### 3. **Best Practices in Verilog Design**
1. **Structured Code**:
   - Maintain a clear structure by separating the module definition, input/output declarations, and functional logic.
   - Use meaningful naming conventions for signals and modules.

2. **Avoiding Latches**:
   - Inadvertent latches can be avoided by ensuring all output paths are covered in combinational logic.
   - All procedural assignments must have values in every conditional branch of control statements.

3. **Simplicity and Clarity**:
   - Use simple and clear logic expressions.
   - Modularize complex designs into smaller, reusable modules.

#### 4. **Common Digital Design Patterns**
1. **Priority Encoder**:
   - Transforms an input vector where several bits might be high, into a binary representation of the highest-priority bit set.
   - Can use a behavioral style with `if-else` or `case` statements to implement priority checking.

2. **State Machines**:
   - Finite State Machines (FSM) control complex sequences of operations.
   - Consist of state definitions, state transitions, and output logic based on current states.

3. **Multiplexers (MUX)**:
   - Selects one of several input signals based on selector bits.
   - Can be implemented using conditional statements or continuous assignment.

#### 5. **Special Considerations**
1. **Synthesis and Simulation**:
   - Ensure that the design is synthesizable by the target hardware (e.g., FPGA, ASIC).
   - Simulation primarily used for functional verification before synthesis.

2. **Resource Utilization**:
   - Optimize designs to minimize hardware resource usage.

3. **Testbenches**:
   - Essential for verifying the functionality of Verilog modules.
   - Include stimulus generation, output monitoring, and self-checking mechanisms.

#### 6. **Debugging and Verification Tools**
1. **Waveform Viewers and Simulators** (e.g., ModelSim, Vivado Simulator):
   - Utilize these tools to visualize signal changes over time.

2. **Assertions and Error Checking**:
   - Implement assertion statements to catch design errors during simulation.

---

This knowledge base serves as a foundation to guide another language model in generating Verilog modules effectively by incorporating fundamental principles, best practices, and common patterns in digital design with Verilog.

Task:
// Build a 4-bit priority encoder. For this problem, if none of the input bits are high 
// (i.e., input is zero), output zero. Note that a 4-bit number has 16 possible combinations.

// Hint: Using hexadecimal (4'hb) or decimal (4'd11) number literals would save typing vs. binary (4'b1011) literals.

// synthesis verilog_input_version verilog_2001
module top_module (
    input [3:0] in,
    output reg [1:0] pos  );

    // Insert your code here

endmodule

