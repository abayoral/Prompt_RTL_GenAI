
# Verilog Design Knowledgebase for Language Models

This knowledgebase encompasses concepts, principles, best practices, and common patterns in Verilog design. It is aimed at enhancing the performance and effectiveness of language models tasked with generating Verilog modules.

### 1. Basic Concepts:
- **Verilog HDL**: A hardware description language used for modeling electronic systems at various levels of abstraction, primarily used in design, verification, and implementation of digital circuits.
- **Modules**: Fundamental building blocks in Verilog, which encapsulate design functionality. Each module can include inputs, outputs, and internal logic.
- **Signals and Variables**: Signals represent wires and storage elements. They can be `wire` (net) type for continuous assignment or `reg` for procedural assignments controlled by always blocks.

### 2. Common Structures:
- **Module Declaration**: Defines interface (ports) and behavior of the hardware module.
- **Instantiation**: Reuse existing modules by creating instances within a higher-level module.
- **Ports**: Module interfaces categorized into inputs, outputs, and bidirectional ports.
- **Parameterization**: Use of parameters to create configurable modules.

### 3. Datatypes:
- **Scalar Datatypes**: Represents single-bit data (`input`, `output`, `wire`, `reg`).
- **Vector Datatypes**: Represents multi-bit data (`input [N:0]`, `output [N:0]`, `integer`, `real`).
- **Arrays and Memories**: Collections of elements, useful for creating memory blocks or large registers.

### 4. Core Principles:
- **Combinational Logic**: Implemented using continuous assignment statements (e.g., `assign`), representing logic without storage elements.
- **Sequential Logic**: Implemented using procedural blocks (`always`, `initial`), representing logic with storage elements (flip-flops, latches).
- **Hierarchy**: Modular design approach where complex systems are built using simpler submodules.

### 5. Best Practices:
- **Readable and Maintainable Code**: Use meaningful module and signal names, follow consistent indentation, and comment your code where necessary.
- **Parameterization**: Utilize parameters for module configurability, allowing the same module to be reused with different configurations.
- **State Machines**: Use state machines for controlling complex sequencing logic.
- **Synchronous Design**: Prefer synchronous reset and clocked logic to enable reliable and predictable behavior.
- **Code Reusability**: Design reusable modules to build scalable and maintainable systems.

### 6. Common Patterns:
- **Adder/Subtractor**: Adder and subtractor functionality can often be combined by using a control signal to toggle between addition and subtraction.
- **Multiplexers (MUX)**: Used for selecting between multiple inputs based on a select signal.
- **Demultiplexers (DEMUX)**: Opposite of multiplexers, used for distributing data from one input to multiple outputs.
- **Shift Registers**: Used for sequentially shifting data in and out.
- **Counters**: Useful for counting events or clock pulses, implemented using flip-flops and combinational logic.
- **State Machines**: Finite State Machines (FSM) for controlling sequential behavior and managing states.
- **Bitwise Operations**: Use of bitwise operators (`&, |, ^, ~`) for performing operations on data at the bit level.

### 7. Bitwise and Logical Operations:
- **Bitwise AND (`&`)**: Performs logical AND on each bit.
- **Bitwise OR (`|`)**: Performs logical OR on each bit.
- **Bitwise XOR (`^`)**: Performs logical exclusive OR on each bit, useful for conditional inversion.
- **Bitwise NOR (`~|`)**: Performs logical NOR.
- **Bitwise NOT (`~`)**: Inverts all bits.
- **Bitwise XNOR (`~^`)**: Performs logical exclusive NOR on each bit.

### 8. Control Structures:
- **Conditional Statements (`if`, `else`, `case`)**: Control the flow of procedural blocks.
- **Loops (`for`, `while`, `repeat`)**: Allow repetitive execution of code segments.

### 9. Timing and Delays:
- **#delay**: Specify delays in assignments to model propagation delays.
- **`@` (event control)**: Trigger statements based on events (edge of a clock or signal).

### 10. Synthesizability:
- Ensure that the code you write is synthesizable and practical to implement in hardware. Avoid using constructs that are not supported by synthesis tools.

---

This knowledgebase should serve as a foundation to inform and guide the generation of Verilog modules. By embedding these principles and best practices, language models can produce high-quality, reliable, and maintainable Verilog designs.

Task:
// Build the adder-subtractor below.
// You are provided with a 16-bit adder module, which you need to instantiate twice:

module add16 ( input[15:0] a, input[15:0] b, input cin, output[15:0] sum, output cout );

// Use a 32-bit wide XOR gate to invert the b input whenever sub is 1. 
// (This can also be viewed as b[31:0] XORed with sub replicated 32 times.). 
// Also connect the sub input to the carry-in of the adder.

// Hint: An XOR gate can also be viewed as a programmable inverter, where one input controls whether the other should be inverted.

module top_module(
    input [31:0] a,
    input [31:0] b,
    input sub,
    output [31:0] sum
);

	// INsert your code here

endmodule