module top_module(
    input a,
    input b,
    input c,
    output out
); 

    // Simplified equation from the Karnaugh map
    assign out = 1;

endmodule