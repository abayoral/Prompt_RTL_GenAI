module top_module(
    output zero
);

    assign zero = 0; // Continuously assign the value 0 to the output 'zero'

endmodule