Please elaborate on the process and code required to create a half adder using Verilog. A half adder is a fundamental arithmetic circuit in digital electronics that adds two single-bit binary numbers (with no carry-in) and outputs two results: a sum bit and a carry-out bit.

Using the provided module template:

```verilog
module top_module( 
    input a, b,
    output cout, sum );
    
    // Insert your code here

endmodule
```

Explain the following elements in your answer:

1. **Purpose of a Half Adder:** What is the primary function of a half adder in digital circuits?
2. **Inputs and Outputs:** Clarify the roles of the inputs `a` and `b`, and the outputs `sum` and `cout`.
3. **Logic and Operations in Half Adder:** Describe the logical operations (such as AND, OR, and XOR) used to determine the values of `sum` and `cout`.
4. **Verilog Implementation:** Guide on how to use Verilog syntax to implement these logical operations properly within the module.

Ensure the explanation is clear enough for someone with basic understanding of digital logic design and Verilog coding standards.