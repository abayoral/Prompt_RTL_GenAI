// you're a senior Digital Design Engineer at a leading hardware design company tasked with developing a critical Verilog module for a next-generation product. The success of this module is pivotal for maintaining my computer hardware company's reputation in the industry.

// Build a combinational circuit with four inputs, in[3:0].

// There are 3 outputs as follows:
// out_and: output of a 4-input AND gate.
// out_or: output of a 4-input OR gate.
// out_xor: output of a 4-input XOR gate.


module top_module( 
    input [3:0] in,
    output out_and,
    output out_or,
    output out_xor
);

// Insert your code here

endmodule