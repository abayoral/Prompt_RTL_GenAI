module top_module( input in, output out );

    // Assign the input signal 'in' to the output signal 'out'
    assign out = in; 

endmodule