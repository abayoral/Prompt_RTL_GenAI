Imagine you are a senior digital design engineer at a leading hardware company, and you’ve been assigned to create a vital Verilog module for an upcoming next-generation computer product. Your task is to develop a D flip-flop circuit that incorporates an asynchronous reset, a design element crucial for the reliable operation of the end product. The module must adhere to strict performance and reliability standards so as to uphold the company’s reputation in the competitive hardware industry.

In this project, you are provided with a module template named "top_module", which includes inputs for the system clock (clk), the data (d), and an asynchronous reset signal (ar), as well as an output (q) representing the flip-flop’s stored state. Your goal is to complete the Verilog code such that it correctly implements the functionality of a D flip-flop with an asynchronous reset. The asynchronous reset must override any other signals and promptly reset the flip-flop output regardless of the clock state. This design will play a pivotal role in the overall performance of the computer hardware product.

The challenge is to write a clear, well-organized, and industry-standard Verilog implementation within the provided module structure, ensuring that all functional requirements—especially the behavior of the asynchronous reset—are accurately met. Note that you are not required to develop any additional features beyond what is specified in this design task.

Remember, no solutions or code should be provided here—only a thorough understanding of the problem and clarification of the design objectives are needed.