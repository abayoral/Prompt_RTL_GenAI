As a senior Digital Design Engineer at a prominent company specializing in hardware design, you have been assigned the crucial task of developing a Verilog module that plays an essential role in a next-generation product. The success of this module is of utmost importance because it significantly impacts your company's standing and reputation in the highly competitive computer hardware industry.

The module you are developing is required to interpret the PS/2 mouse protocol, which organizes its communication into messages that are precisely three bytes long. One challenging aspect of working with this protocol is the nature of the byte stream; it does not clearly indicate where individual messages begin and end. The only distinctive feature that signals the start of a new message is the first byte, which has bit[3] set to 1. In contrast, the bits[3] of the subsequent two bytes may either be 1 or 0, depending on the data being transmitted.

With this understanding, your task is to design a finite state machine (FSM) that effectively searches for the boundaries of these messages within an incoming byte stream. The proposed algorithm suggests that the FSM should actively discard any incoming bytes until it encounters a byte where bit[3] equals 1. This byte is assumed to be the first part of a new message, and the FSM needs to signal the completion of a message only after receiving all three bytes, which would then result in asserting the `done` signal.

As part of your design specifications, it is essential that the FSM indicates that a message has been completely received during the clock cycle following the reception of the third byte. While the input `in[7:0]` represents a single byte, the FSM must primarily utilize only the value of bit[3] from this byte for its state transitions. You anticipate needing approximately four states to manage this process effectively. This number is necessary because at least one of those states must be responsible for asserting the `done` signal, and this signal should only be active for one clock cycle corresponding to each received message.

With these requirements in mind, how would you approach the design and implementation of this FSM in your Verilog module? What considerations might influence the state transition logic, the defining of the states within the FSM, and the output logic necessary for signaling the completion of each message? Additionally, how would you organize the sequential elements of the FSM to respond appropriately to the incoming byte stream while ensuring that the reset functionality operates as intended?